module top(
  input logic [23:0] x_i, y_i,
/* verilator lint_off UNUSED */
  input logic clk_i,
  output logic [23:0] z_o
);

modular_mul dut(.*);

endmodule: top
